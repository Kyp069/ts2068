//-------------------------------------------------------------------------------------------------
module dprs
//-------------------------------------------------------------------------------------------------
#
(
	parameter KB = 0
)
(
	input  wire                      clock1,
	input  wire[$clog2(KB*1024)-1:0] a1,
	output reg [                7:0] q1,
	input  wire                      clock2,
	input  wire[$clog2(KB*1024)-1:0] a2,
	input  wire[                7:0] d2,
	input  wire                      w2
);
//-------------------------------------------------------------------------------------------------

reg[7:0] mem[0:(KB*1024)-1];

wire w1 = 1'b0;
wire[7:0] d1 = 8'hFF;

always @(posedge clock1) if(w1) begin q1 <= d1; mem[a1] <= d1; end else q1 <= mem[a1];
always @(posedge clock2) if(w2) mem[a2] <= d2;

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------
module dprf
//-------------------------------------------------------------------------------------------------
#
(
	parameter KB = 0
)
(
	input  wire                      clock1,
	input  wire[$clog2(KB*1024)-1:0] a1,
	output reg [                7:0] q1,
	input  wire                      clock2,
	input  wire[$clog2(KB*1024)-1:0] a2,
	input  wire[                7:0] d2,
	output reg [                7:0] q2,
	input  wire                      w2
);
//-------------------------------------------------------------------------------------------------

reg[7:0] mem[0:(KB*1024)-1];

wire w1 = 1'b0;
wire[7:0] d1 = 8'hFF;

always @(posedge clock1) if(w1) begin q1 <= d1; mem[a1] <= d1; end else q1 <= mem[a1];
always @(posedge clock2) if(w2) begin q2 <= d2; mem[a2] <= d2; end else q2 <= mem[a2];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------
module dprfm
//-------------------------------------------------------------------------------------------------
#
(
	parameter KB = 0,
	parameter FN = ""
)
(
	input  wire                      clock1,
	input  wire[$clog2(KB*1024)-1:0] a1,
	output reg [                7:0] q1,
	input  wire                      clock2,
	input  wire[$clog2(KB*1024)-1:0] a2,
	input  wire[                7:0] d2,
	output reg [                7:0] q2,
	input  wire                      w2
);
//-------------------------------------------------------------------------------------------------

(* ram_init_file = FN *) reg[7:0] mem[0:(KB*1024)-1];

wire w1 = 1'b0;
wire[7:0] d1 = 8'hFF;

always @(posedge clock1) if(w1) begin q1 <= d1; mem[a1] <= d1; end else q1 <= mem[a1];
always @(posedge clock2) if(w2) begin q2 <= d2; mem[a2] <= d2; end else q2 <= mem[a2];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------

// reg[7:0] mem[0:(KB*1024)-1] /* synthesis ram_init_file = FN */;
// initial if(FN != "") $readmemh(FN, mem);
